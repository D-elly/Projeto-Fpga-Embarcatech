module eff_1( 

);

endmodule